interface flip_flop;
  
  logic clk;
  
  logic rst_n;
  
  logic data;
  
  logic q;
  
  logic q_bar;
  
endinterface
